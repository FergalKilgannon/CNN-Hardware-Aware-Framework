`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company:       	UCD School of Electrical and Electronic Engineering
// Student:   		Fergal Kilgannon
// Student num:	  	19315126
// Project:       	CNN Hardware-Software Codesign
// Description:   	Digital Multiply-and-Accumulate module testbench
// Last edited:   	26th December 2023
//////////////////////////////////////////////////////////////////////////////////

module TBlinearMAC;

	reg clock, reset, enable;
	reg [7:0] data_in, weight_in;
	
	wire [16:0] result;
  
  // Integer variable to count errors
	integer error_count;
	
// Instantiate top level module
	digital_MAC uut (
		.clock(clock),
		.data_in(data_in),
		.weight_in(weight_in),
		.reset(reset),
      	.enable(enable),
		.data_out(result)
	);

// Generate clock signal at 250 MHz
	initial 
		begin
			clock = 1'b0;  // clock starts at 0
			forever
				#4 clock = ~clock;	// invert clock every 4 ns
		end
		
	initial 
      begin
				reset = 1'b0;
				data_in = 15'b0;
				weight_in = 15'b0;
        enable = 1'b0;
        error_count = 0;	// initialise error counter
        
        #4;
				reset = 1'b1;
      	@ (negedge clock);
      	@ (negedge clock) reset = 1'b0;
		
		// Start of custom
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd84, -15'd82);
        #4;
        CHECK_ACCUM(15'd-6888);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd84, -15'd91);
        #4;
        MULT(15'd222, -15'd82);
        #4;
        CHECK_ACCUM(15'd-25848);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd84, -15'd9);
        #4;
        MULT(15'd222, -15'd91);
        #4;
        MULT(15'd67, -15'd82);
        #4;
        CHECK_ACCUM(15'd-26452);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd84, 15'd102);
        #4;
        MULT(15'd222, -15'd9);
        #4;
        MULT(15'd67, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd473);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd84, -15'd38);
        #4;
        MULT(15'd222, 15'd102);
        #4;
        MULT(15'd67, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd18849);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd222, -15'd38);
        #4;
        MULT(15'd67, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1602);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd67, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2546);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd84, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd185, -15'd82);
        #4;
        CHECK_ACCUM(15'd286);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd84, 15'd197);
        #4;
        MULT(15'd222, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd185, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd19733);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd84, 15'd169);
        #4;
        MULT(15'd222, 15'd197);
        #4;
        MULT(15'd67, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd185, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd114, -15'd82);
        #4;
        CHECK_ACCUM(15'd36131);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd84, 15'd105);
        #4;
        MULT(15'd222, 15'd169);
        #4;
        MULT(15'd67, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd185, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd114, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd65747);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd84, 15'd60);
        #4;
        MULT(15'd222, 15'd105);
        #4;
        MULT(15'd67, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd185, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd114, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd57525);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd222, 15'd60);
        #4;
        MULT(15'd67, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd114, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd22331);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd67, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd114, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-312);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd84, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd185, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd159, -15'd82);
        #4;
        CHECK_ACCUM(15'd22598);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd84, 15'd55);
        #4;
        MULT(15'd222, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd185, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd159, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd56722);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd84, 15'd55);
        #4;
        MULT(15'd222, 15'd55);
        #4;
        MULT(15'd67, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd185, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd114, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd159, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd72, -15'd82);
        #4;
        CHECK_ACCUM(15'd89933);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd84, 15'd7);
        #4;
        MULT(15'd222, 15'd55);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd185, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd114, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd159, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd72, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd108672);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd84, -15'd19);
        #4;
        MULT(15'd222, 15'd7);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd185, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd114, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd159, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd72, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd79897);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd222, -15'd19);
        #4;
        MULT(15'd67, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd114, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd72, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd21153);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd67, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd114, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd72, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd2831);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd84, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd185, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd159, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd151, -15'd82);
        #4;
        CHECK_ACCUM(15'd17365);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd84, -15'd61);
        #4;
        MULT(15'd222, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd185, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd159, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd151, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd45375);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd84, -15'd100);
        #4;
        MULT(15'd222, -15'd61);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd185, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd114, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd159, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd72, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd151, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd114, -15'd82);
        #4;
        CHECK_ACCUM(15'd58293);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd84, -15'd92);
        #4;
        MULT(15'd222, -15'd100);
        #4;
        MULT(15'd67, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd185, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd114, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd159, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd72, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd151, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd114, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd64067);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd84, -15'd8);
        #4;
        MULT(15'd222, -15'd92);
        #4;
        MULT(15'd67, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd185, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd114, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd159, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd72, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd151, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd114, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd44259);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd222, -15'd8);
        #4;
        MULT(15'd67, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd114, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd72, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd114, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd12808);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd67, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd114, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd72, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd114, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2714);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd84, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd185, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd159, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd151, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd60, -15'd82);
        #4;
        CHECK_ACCUM(15'd10321);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd84, -15'd3);
        #4;
        MULT(15'd222, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd185, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd159, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd151, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd60, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd19553);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd84, -15'd144);
        #4;
        MULT(15'd222, -15'd3);
        #4;
        MULT(15'd67, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd185, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd114, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd159, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd72, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd151, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd114, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd60, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd163, -15'd82);
        #4;
        CHECK_ACCUM(15'd25634);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd84, -15'd120);
        #4;
        MULT(15'd222, -15'd144);
        #4;
        MULT(15'd67, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd185, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd114, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd159, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd72, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd151, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd114, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd60, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd163, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2340);
        #4;
        MULT(15'd84, -15'd36);
        #4;
        MULT(15'd222, -15'd120);
        #4;
        MULT(15'd67, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd185, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd114, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd159, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd72, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd151, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd114, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd60, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd163, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd4314);
        #4;
        MULT(15'd222, -15'd36);
        #4;
        MULT(15'd67, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd114, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd72, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd114, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd163, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd1310);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd114, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd72, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd114, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd163, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-4046);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd61, -15'd82);
        #4;
        CHECK_ACCUM(15'd-5002);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd61, -15'd91);
        #4;
        MULT(15'd121, -15'd82);
        #4;
        CHECK_ACCUM(15'd-15473);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd61, -15'd9);
        #4;
        MULT(15'd121, -15'd91);
        #4;
        MULT(15'd121, -15'd82);
        #4;
        CHECK_ACCUM(15'd-21482);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd185, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd159, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd151, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd60, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd36, -15'd82);
        #4;
        CHECK_ACCUM(15'd-14377);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd185, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd159, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd151, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd60, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd36, -15'd91);
        #4;
        MULT(15'd241, -15'd82);
        #4;
        CHECK_ACCUM(15'd2327);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd185, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd114, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd159, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd72, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd151, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd114, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd60, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd163, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd36, -15'd9);
        #4;
        MULT(15'd241, -15'd91);
        #4;
        MULT(15'd227, -15'd82);
        #4;
        CHECK_ACCUM(15'd270);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd185, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd114, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd159, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd72, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd151, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd114, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd60, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd163, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd36, 15'd102);
        #4;
        MULT(15'd241, -15'd9);
        #4;
        MULT(15'd227, -15'd91);
        #4;
        MULT(15'd17, -15'd82);
        #4;
        CHECK_ACCUM(15'd-21452);
        #4;
        MULT(15'd185, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd114, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd159, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd72, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd151, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd114, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd60, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd163, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd36, -15'd38);
        #4;
        MULT(15'd241, 15'd102);
        #4;
        MULT(15'd227, -15'd9);
        #4;
        MULT(15'd17, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2776);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd114, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd72, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd114, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd163, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd241, -15'd38);
        #4;
        MULT(15'd227, 15'd102);
        #4;
        MULT(15'd17, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd10690);
        #4;
        MULT(15'd114, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd72, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd114, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd163, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd227, -15'd38);
        #4;
        MULT(15'd17, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-3958);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd17, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-646);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd31, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2542);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd31, -15'd91);
        #4;
        MULT(15'd133, -15'd82);
        #4;
        CHECK_ACCUM(15'd-13727);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd61, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd31, -15'd9);
        #4;
        MULT(15'd133, -15'd91);
        #4;
        MULT(15'd242, -15'd82);
        #4;
        CHECK_ACCUM(15'd-21002);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd61, 15'd197);
        #4;
        MULT(15'd121, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd31, 15'd102);
        #4;
        MULT(15'd133, -15'd9);
        #4;
        MULT(15'd242, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd-6604);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd61, 15'd169);
        #4;
        MULT(15'd121, 15'd197);
        #4;
        MULT(15'd121, 15'd184);
        #4;
        MULT(15'd31, -15'd38);
        #4;
        MULT(15'd133, 15'd102);
        #4;
        MULT(15'd242, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd22678);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd159, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd151, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd60, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd36, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-14526);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd159, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd151, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd60, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd36, 15'd197);
        #4;
        MULT(15'd241, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2430);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd159, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd72, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd151, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd114, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd60, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd163, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd36, 15'd169);
        #4;
        MULT(15'd241, 15'd197);
        #4;
        MULT(15'd227, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd10862);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd159, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd72, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd151, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd114, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd60, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd163, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd36, 15'd105);
        #4;
        MULT(15'd241, 15'd169);
        #4;
        MULT(15'd227, 15'd197);
        #4;
        MULT(15'd17, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd66, -15'd82);
        #4;
        CHECK_ACCUM(15'd-16715);
        #4;
        MULT(15'd159, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd72, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd151, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd114, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd60, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd163, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd36, 15'd60);
        #4;
        MULT(15'd241, 15'd105);
        #4;
        MULT(15'd227, 15'd169);
        #4;
        MULT(15'd17, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd66, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd8136);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd72, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd114, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd163, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd241, 15'd60);
        #4;
        MULT(15'd227, 15'd105);
        #4;
        MULT(15'd17, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd66, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd24969);
        #4;
        MULT(15'd72, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd114, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd163, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd227, 15'd60);
        #4;
        MULT(15'd17, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd66, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd5884);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd17, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd66, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1488);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd3, -15'd82);
        #4;
        CHECK_ACCUM(15'd-246);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd3, -15'd91);
        #4;
        MULT(15'd38, -15'd82);
        #4;
        CHECK_ACCUM(15'd-3389);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd31, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd3, -15'd9);
        #4;
        MULT(15'd38, -15'd91);
        #4;
        MULT(15'd224, -15'd82);
        #4;
        CHECK_ACCUM(15'd-16149);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd31, 15'd197);
        #4;
        MULT(15'd133, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd3, 15'd102);
        #4;
        MULT(15'd38, -15'd9);
        #4;
        MULT(15'd224, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd-10669);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd61, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd31, 15'd169);
        #4;
        MULT(15'd133, 15'd197);
        #4;
        MULT(15'd242, 15'd184);
        #4;
        MULT(15'd3, -15'd38);
        #4;
        MULT(15'd38, 15'd102);
        #4;
        MULT(15'd224, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd34931);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd61, 15'd55);
        #4;
        MULT(15'd121, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd31, 15'd105);
        #4;
        MULT(15'd133, 15'd169);
        #4;
        MULT(15'd242, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd38, -15'd38);
        #4;
        MULT(15'd224, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd100972);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd61, 15'd55);
        #4;
        MULT(15'd121, 15'd55);
        #4;
        MULT(15'd121, 15'd19);
        #4;
        MULT(15'd31, 15'd60);
        #4;
        MULT(15'd133, 15'd105);
        #4;
        MULT(15'd242, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd224, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd207, -15'd82);
        #4;
        CHECK_ACCUM(15'd140828);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd151, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd60, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd36, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-17482);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd151, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd60, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd36, 15'd55);
        #4;
        MULT(15'd241, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-13426);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd151, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd114, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd60, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd163, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd36, 15'd55);
        #4;
        MULT(15'd241, 15'd55);
        #4;
        MULT(15'd227, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd225, -15'd82);
        #4;
        CHECK_ACCUM(15'd6870);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd151, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd114, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd60, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd163, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd36, 15'd7);
        #4;
        MULT(15'd241, 15'd55);
        #4;
        MULT(15'd227, 15'd55);
        #4;
        MULT(15'd17, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd66, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd225, -15'd91);
        #4;
        MULT(15'd14, -15'd82);
        #4;
        CHECK_ACCUM(15'd2653);
        #4;
        MULT(15'd151, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd114, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd60, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd163, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd36, -15'd19);
        #4;
        MULT(15'd241, 15'd7);
        #4;
        MULT(15'd227, 15'd55);
        #4;
        MULT(15'd17, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd66, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd225, -15'd9);
        #4;
        MULT(15'd14, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd15558);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd114, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd163, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd241, -15'd19);
        #4;
        MULT(15'd227, 15'd7);
        #4;
        MULT(15'd17, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd66, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd225, 15'd102);
        #4;
        MULT(15'd14, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd23097);
        #4;
        MULT(15'd114, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd163, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd227, -15'd19);
        #4;
        MULT(15'd17, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd66, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd225, -15'd38);
        #4;
        MULT(15'd14, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd5446);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd17, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd66, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd14, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd3105);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd19, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1558);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd3, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd19, -15'd91);
        #4;
        MULT(15'd203, -15'd82);
        #4;
        CHECK_ACCUM(15'd-17823);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd3, 15'd197);
        #4;
        MULT(15'd38, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd19, -15'd9);
        #4;
        MULT(15'd203, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd-31889);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd31, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd3, 15'd169);
        #4;
        MULT(15'd38, 15'd197);
        #4;
        MULT(15'd224, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd19, 15'd102);
        #4;
        MULT(15'd203, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd5967);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd31, 15'd55);
        #4;
        MULT(15'd133, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd3, 15'd105);
        #4;
        MULT(15'd38, 15'd169);
        #4;
        MULT(15'd224, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd19, -15'd38);
        #4;
        MULT(15'd203, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd75589);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd61, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd31, 15'd55);
        #4;
        MULT(15'd133, 15'd55);
        #4;
        MULT(15'd242, 15'd19);
        #4;
        MULT(15'd3, 15'd60);
        #4;
        MULT(15'd38, 15'd105);
        #4;
        MULT(15'd224, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd203, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd122188);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd61, -15'd61);
        #4;
        MULT(15'd121, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd31, 15'd7);
        #4;
        MULT(15'd133, 15'd55);
        #4;
        MULT(15'd242, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd38, 15'd60);
        #4;
        MULT(15'd224, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd219, -15'd82);
        #4;
        CHECK_ACCUM(15'd155989);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd61, -15'd100);
        #4;
        MULT(15'd121, -15'd61);
        #4;
        MULT(15'd121, -15'd36);
        #4;
        MULT(15'd31, -15'd19);
        #4;
        MULT(15'd133, 15'd7);
        #4;
        MULT(15'd242, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd224, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd207, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd219, -15'd91);
        #4;
        MULT(15'd18, -15'd82);
        #4;
        CHECK_ACCUM(15'd178338);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd60, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd36, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-7656);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd60, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd36, -15'd61);
        #4;
        MULT(15'd241, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-14018);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd60, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd163, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd36, -15'd100);
        #4;
        MULT(15'd241, -15'd61);
        #4;
        MULT(15'd227, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd225, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd4123);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd60, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd163, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd36, -15'd92);
        #4;
        MULT(15'd241, -15'd100);
        #4;
        MULT(15'd227, -15'd61);
        #4;
        MULT(15'd17, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd66, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd225, 15'd197);
        #4;
        MULT(15'd14, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd67, -15'd82);
        #4;
        CHECK_ACCUM(15'd-10049);
        #4;
        MULT(15'd60, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd163, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd36, -15'd8);
        #4;
        MULT(15'd241, -15'd92);
        #4;
        MULT(15'd227, -15'd100);
        #4;
        MULT(15'd17, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd66, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd225, 15'd169);
        #4;
        MULT(15'd14, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd67, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-9937);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd163, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd241, -15'd8);
        #4;
        MULT(15'd227, -15'd92);
        #4;
        MULT(15'd17, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd66, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd225, 15'd105);
        #4;
        MULT(15'd14, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd67, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd4082);
        #4;
        MULT(15'd163, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd227, -15'd8);
        #4;
        MULT(15'd17, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd66, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd225, 15'd60);
        #4;
        MULT(15'd14, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd67, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1460);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd17, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd66, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd14, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd67, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-3096);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd75, -15'd82);
        #4;
        CHECK_ACCUM(15'd-6150);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd19, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd75, -15'd91);
        #4;
        MULT(15'd221, -15'd82);
        #4;
        CHECK_ACCUM(15'd-21451);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd3, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd19, 15'd197);
        #4;
        MULT(15'd203, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd75, -15'd9);
        #4;
        MULT(15'd221, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd-462);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd3, 15'd55);
        #4;
        MULT(15'd38, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd19, 15'd169);
        #4;
        MULT(15'd203, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd75, 15'd102);
        #4;
        MULT(15'd221, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd52544);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd31, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd3, 15'd55);
        #4;
        MULT(15'd38, 15'd55);
        #4;
        MULT(15'd224, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd19, 15'd105);
        #4;
        MULT(15'd203, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd75, -15'd38);
        #4;
        MULT(15'd221, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd115, -15'd82);
        #4;
        CHECK_ACCUM(15'd123333);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd31, -15'd61);
        #4;
        MULT(15'd133, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd3, 15'd7);
        #4;
        MULT(15'd38, 15'd55);
        #4;
        MULT(15'd224, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd19, 15'd60);
        #4;
        MULT(15'd203, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd221, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd115, -15'd91);
        #4;
        MULT(15'd52, -15'd82);
        #4;
        CHECK_ACCUM(15'd175228);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd61, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd31, -15'd100);
        #4;
        MULT(15'd133, -15'd61);
        #4;
        MULT(15'd242, -15'd36);
        #4;
        MULT(15'd3, -15'd19);
        #4;
        MULT(15'd38, 15'd7);
        #4;
        MULT(15'd224, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd203, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd115, -15'd9);
        #4;
        MULT(15'd52, -15'd91);
        #4;
        MULT(15'd52, -15'd82);
        #4;
        CHECK_ACCUM(15'd189709);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd61, -15'd3);
        #4;
        MULT(15'd121, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd31, -15'd92);
        #4;
        MULT(15'd133, -15'd100);
        #4;
        MULT(15'd242, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd38, -15'd19);
        #4;
        MULT(15'd224, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd219, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd115, 15'd102);
        #4;
        MULT(15'd52, -15'd9);
        #4;
        MULT(15'd52, -15'd91);
        #4;
        MULT(15'd40, -15'd82);
        #4;
        CHECK_ACCUM(15'd149313);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd61, -15'd144);
        #4;
        MULT(15'd121, -15'd3);
        #4;
        MULT(15'd121, -15'd106);
        #4;
        MULT(15'd31, -15'd8);
        #4;
        MULT(15'd133, -15'd92);
        #4;
        MULT(15'd242, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd224, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd207, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd219, 15'd197);
        #4;
        MULT(15'd18, 15'd184);
        #4;
        MULT(15'd115, -15'd38);
        #4;
        MULT(15'd52, 15'd102);
        #4;
        MULT(15'd52, -15'd9);
        #4;
        MULT(15'd40, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd74217);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd36, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-3816);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd36, -15'd3);
        #4;
        MULT(15'd241, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-8824);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd36, -15'd144);
        #4;
        MULT(15'd241, -15'd3);
        #4;
        MULT(15'd227, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd225, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd10870);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd36, -15'd120);
        #4;
        MULT(15'd241, -15'd144);
        #4;
        MULT(15'd227, -15'd3);
        #4;
        MULT(15'd17, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd66, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd225, 15'd55);
        #4;
        MULT(15'd14, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd67, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd67, -15'd82);
        #4;
        CHECK_ACCUM(15'd9792);
        #4;
        MULT(15'd36, -15'd36);
        #4;
        MULT(15'd241, -15'd120);
        #4;
        MULT(15'd227, -15'd144);
        #4;
        MULT(15'd17, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd66, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd225, 15'd55);
        #4;
        MULT(15'd14, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd67, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd67, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-7338);
        #4;
        MULT(15'd241, -15'd36);
        #4;
        MULT(15'd227, -15'd120);
        #4;
        MULT(15'd17, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd66, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd225, 15'd7);
        #4;
        MULT(15'd14, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd67, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd67, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-3679);
        #4;
        MULT(15'd227, -15'd36);
        #4;
        MULT(15'd17, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd66, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd225, -15'd19);
        #4;
        MULT(15'd14, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd67, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd67, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-3036);
        #4;
        MULT(15'd17, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd66, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd14, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd67, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd67, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd68);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd9, -15'd82);
        #4;
        CHECK_ACCUM(15'd-738);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd9, -15'd91);
        #4;
        MULT(15'd126, -15'd82);
        #4;
        CHECK_ACCUM(15'd-11151);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd75, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd9, -15'd9);
        #4;
        MULT(15'd126, -15'd91);
        #4;
        MULT(15'd251, -15'd82);
        #4;
        CHECK_ACCUM(15'd-18329);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd19, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd75, 15'd197);
        #4;
        MULT(15'd221, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd9, 15'd102);
        #4;
        MULT(15'd126, -15'd9);
        #4;
        MULT(15'd251, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd11915);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd3, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd19, 15'd55);
        #4;
        MULT(15'd203, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd75, 15'd169);
        #4;
        MULT(15'd221, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd9, -15'd38);
        #4;
        MULT(15'd126, 15'd102);
        #4;
        MULT(15'd251, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd219, -15'd82);
        #4;
        CHECK_ACCUM(15'd76921);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd3, -15'd61);
        #4;
        MULT(15'd38, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd19, 15'd55);
        #4;
        MULT(15'd203, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd75, 15'd105);
        #4;
        MULT(15'd221, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd126, -15'd38);
        #4;
        MULT(15'd251, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd219, -15'd91);
        #4;
        MULT(15'd77, -15'd82);
        #4;
        CHECK_ACCUM(15'd149768);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd31, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd3, -15'd100);
        #4;
        MULT(15'd38, -15'd61);
        #4;
        MULT(15'd224, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd19, 15'd7);
        #4;
        MULT(15'd203, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd75, 15'd60);
        #4;
        MULT(15'd221, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd115, 15'd184);
        #4;
        MULT(15'd251, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd219, -15'd9);
        #4;
        MULT(15'd77, -15'd91);
        #4;
        MULT(15'd1, -15'd82);
        #4;
        CHECK_ACCUM(15'd165265);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd31, -15'd3);
        #4;
        MULT(15'd133, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd3, -15'd92);
        #4;
        MULT(15'd38, -15'd100);
        #4;
        MULT(15'd224, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd19, -15'd19);
        #4;
        MULT(15'd203, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd221, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd115, 15'd197);
        #4;
        MULT(15'd52, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd219, 15'd102);
        #4;
        MULT(15'd77, -15'd9);
        #4;
        MULT(15'd1, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd119732);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd31, -15'd144);
        #4;
        MULT(15'd133, -15'd3);
        #4;
        MULT(15'd242, -15'd106);
        #4;
        MULT(15'd3, -15'd8);
        #4;
        MULT(15'd38, -15'd92);
        #4;
        MULT(15'd224, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd203, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd115, 15'd169);
        #4;
        MULT(15'd52, 15'd197);
        #4;
        MULT(15'd52, 15'd184);
        #4;
        MULT(15'd219, -15'd38);
        #4;
        MULT(15'd77, 15'd102);
        #4;
        MULT(15'd1, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd30294);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd31, -15'd120);
        #4;
        MULT(15'd133, -15'd144);
        #4;
        MULT(15'd242, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd38, -15'd8);
        #4;
        MULT(15'd224, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd219, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd115, 15'd105);
        #4;
        MULT(15'd52, 15'd169);
        #4;
        MULT(15'd52, 15'd197);
        #4;
        MULT(15'd40, 15'd184);
        #4;
        MULT(15'd77, -15'd38);
        #4;
        MULT(15'd1, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-41536);
        #4;
        MULT(15'd31, -15'd36);
        #4;
        MULT(15'd133, -15'd120);
        #4;
        MULT(15'd242, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd224, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd207, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd219, 15'd55);
        #4;
        MULT(15'd18, 15'd19);
        #4;
        MULT(15'd115, 15'd60);
        #4;
        MULT(15'd52, 15'd105);
        #4;
        MULT(15'd52, 15'd169);
        #4;
        MULT(15'd40, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd1, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-100817);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-4158);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd225, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd14916);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd66, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd225, -15'd61);
        #4;
        MULT(15'd14, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd67, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd67, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd67, -15'd82);
        #4;
        CHECK_ACCUM(15'd21272);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd66, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd225, -15'd100);
        #4;
        MULT(15'd14, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd67, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd67, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd5665);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd66, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd225, -15'd92);
        #4;
        MULT(15'd14, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd67, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd67, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1441);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd66, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd225, -15'd8);
        #4;
        MULT(15'd14, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd67, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd67, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd67, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-5052);
        #4;
        MULT(15'd66, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd14, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd67, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd67, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd67, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd59, -15'd82);
        #4;
        CHECK_ACCUM(15'd-7125);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd59, -15'd91);
        #4;
        MULT(15'd133, -15'd82);
        #4;
        CHECK_ACCUM(15'd-16275);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd9, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd59, -15'd9);
        #4;
        MULT(15'd133, -15'd91);
        #4;
        MULT(15'd205, -15'd82);
        #4;
        CHECK_ACCUM(15'd-27788);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd9, 15'd197);
        #4;
        MULT(15'd126, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd59, 15'd102);
        #4;
        MULT(15'd133, -15'd9);
        #4;
        MULT(15'd205, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd-9705);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd75, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd9, 15'd169);
        #4;
        MULT(15'd126, 15'd197);
        #4;
        MULT(15'd251, 15'd184);
        #4;
        MULT(15'd59, -15'd38);
        #4;
        MULT(15'd133, 15'd102);
        #4;
        MULT(15'd205, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd240, -15'd82);
        #4;
        CHECK_ACCUM(15'd40637);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd19, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd75, 15'd55);
        #4;
        MULT(15'd221, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd9, 15'd105);
        #4;
        MULT(15'd126, 15'd169);
        #4;
        MULT(15'd251, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd133, -15'd38);
        #4;
        MULT(15'd205, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd240, -15'd91);
        #4;
        MULT(15'd166, -15'd82);
        #4;
        CHECK_ACCUM(15'd104180);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd3, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd19, -15'd61);
        #4;
        MULT(15'd203, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd75, 15'd55);
        #4;
        MULT(15'd221, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd9, 15'd60);
        #4;
        MULT(15'd126, 15'd105);
        #4;
        MULT(15'd251, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd219, 15'd184);
        #4;
        MULT(15'd205, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd240, -15'd9);
        #4;
        MULT(15'd166, -15'd91);
        #4;
        MULT(15'd35, -15'd82);
        #4;
        CHECK_ACCUM(15'd156826);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd3, -15'd3);
        #4;
        MULT(15'd38, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd19, -15'd100);
        #4;
        MULT(15'd203, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd75, 15'd7);
        #4;
        MULT(15'd221, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd126, 15'd60);
        #4;
        MULT(15'd251, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd219, 15'd197);
        #4;
        MULT(15'd77, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd240, 15'd102);
        #4;
        MULT(15'd166, -15'd9);
        #4;
        MULT(15'd35, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd148313);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd3, -15'd144);
        #4;
        MULT(15'd38, -15'd3);
        #4;
        MULT(15'd224, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd19, -15'd92);
        #4;
        MULT(15'd203, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd75, -15'd19);
        #4;
        MULT(15'd221, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd115, 15'd19);
        #4;
        MULT(15'd251, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd219, 15'd169);
        #4;
        MULT(15'd77, 15'd197);
        #4;
        MULT(15'd1, 15'd184);
        #4;
        MULT(15'd240, -15'd38);
        #4;
        MULT(15'd166, 15'd102);
        #4;
        MULT(15'd35, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd60862);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd3, -15'd120);
        #4;
        MULT(15'd38, -15'd144);
        #4;
        MULT(15'd224, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd19, -15'd8);
        #4;
        MULT(15'd203, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd221, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd115, 15'd55);
        #4;
        MULT(15'd52, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd219, 15'd105);
        #4;
        MULT(15'd77, 15'd169);
        #4;
        MULT(15'd1, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd166, -15'd38);
        #4;
        MULT(15'd35, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-34725);
        #4;
        MULT(15'd3, -15'd36);
        #4;
        MULT(15'd38, -15'd120);
        #4;
        MULT(15'd224, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd203, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd115, 15'd55);
        #4;
        MULT(15'd52, 15'd55);
        #4;
        MULT(15'd52, 15'd19);
        #4;
        MULT(15'd219, 15'd60);
        #4;
        MULT(15'd77, 15'd105);
        #4;
        MULT(15'd1, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd35, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-112451);
        #4;
        MULT(15'd38, -15'd36);
        #4;
        MULT(15'd224, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd219, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd115, 15'd7);
        #4;
        MULT(15'd52, 15'd55);
        #4;
        MULT(15'd52, 15'd55);
        #4;
        MULT(15'd40, 15'd19);
        #4;
        MULT(15'd77, 15'd60);
        #4;
        MULT(15'd1, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-159504);
        #4;
        MULT(15'd224, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd207, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd219, -15'd61);
        #4;
        MULT(15'd18, -15'd36);
        #4;
        MULT(15'd115, -15'd19);
        #4;
        MULT(15'd52, 15'd7);
        #4;
        MULT(15'd52, 15'd55);
        #4;
        MULT(15'd40, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd1, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-159332);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-4158);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd225, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd250, -15'd82);
        #4;
        CHECK_ACCUM(15'd17274);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd225, -15'd3);
        #4;
        MULT(15'd14, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd67, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd67, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd250, -15'd91);
        #4;
        MULT(15'd59, -15'd82);
        #4;
        CHECK_ACCUM(15'd24214);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd225, -15'd144);
        #4;
        MULT(15'd14, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd67, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd67, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd250, -15'd9);
        #4;
        MULT(15'd59, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd4628);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd225, -15'd120);
        #4;
        MULT(15'd14, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd67, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd67, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd250, 15'd102);
        #4;
        MULT(15'd59, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd22, -15'd82);
        #4;
        CHECK_ACCUM(15'd-581);
        #4;
        MULT(15'd225, -15'd36);
        #4;
        MULT(15'd14, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd67, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd67, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd67, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd250, -15'd38);
        #4;
        MULT(15'd59, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd22, -15'd91);
        #4;
        MULT(15'd129, -15'd82);
        #4;
        CHECK_ACCUM(15'd-16120);
        #4;
        MULT(15'd14, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd67, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd67, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd67, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd59, 15'd184);
        #4;
        MULT(15'd59, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd22, -15'd9);
        #4;
        MULT(15'd129, -15'd91);
        #4;
        MULT(15'd249, -15'd82);
        #4;
        CHECK_ACCUM(15'd-22034);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd59, 15'd197);
        #4;
        MULT(15'd133, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd22, 15'd102);
        #4;
        MULT(15'd129, -15'd9);
        #4;
        MULT(15'd249, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd-6309);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd9, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd59, 15'd169);
        #4;
        MULT(15'd133, 15'd197);
        #4;
        MULT(15'd205, 15'd184);
        #4;
        MULT(15'd22, -15'd38);
        #4;
        MULT(15'd129, 15'd102);
        #4;
        MULT(15'd249, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd248, -15'd82);
        #4;
        CHECK_ACCUM(15'd40694);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd9, 15'd55);
        #4;
        MULT(15'd126, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd59, 15'd105);
        #4;
        MULT(15'd133, 15'd169);
        #4;
        MULT(15'd205, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd129, -15'd38);
        #4;
        MULT(15'd249, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd248, -15'd91);
        #4;
        MULT(15'd182, -15'd82);
        #4;
        CHECK_ACCUM(15'd99400);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd75, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd9, 15'd55);
        #4;
        MULT(15'd126, 15'd55);
        #4;
        MULT(15'd251, 15'd19);
        #4;
        MULT(15'd59, 15'd60);
        #4;
        MULT(15'd133, 15'd105);
        #4;
        MULT(15'd205, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd240, 15'd184);
        #4;
        MULT(15'd249, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd248, -15'd9);
        #4;
        MULT(15'd182, -15'd91);
        #4;
        MULT(15'd57, -15'd82);
        #4;
        CHECK_ACCUM(15'd148820);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd19, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd75, -15'd61);
        #4;
        MULT(15'd221, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd9, 15'd7);
        #4;
        MULT(15'd126, 15'd55);
        #4;
        MULT(15'd251, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd133, 15'd60);
        #4;
        MULT(15'd205, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd240, 15'd197);
        #4;
        MULT(15'd166, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd248, 15'd102);
        #4;
        MULT(15'd182, -15'd9);
        #4;
        MULT(15'd57, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd170153);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd19, -15'd3);
        #4;
        MULT(15'd203, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd75, -15'd100);
        #4;
        MULT(15'd221, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd9, -15'd19);
        #4;
        MULT(15'd126, 15'd7);
        #4;
        MULT(15'd251, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd219, 15'd19);
        #4;
        MULT(15'd205, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd240, 15'd169);
        #4;
        MULT(15'd166, 15'd197);
        #4;
        MULT(15'd35, 15'd184);
        #4;
        MULT(15'd248, -15'd38);
        #4;
        MULT(15'd182, 15'd102);
        #4;
        MULT(15'd57, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd108246);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd19, -15'd144);
        #4;
        MULT(15'd203, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd75, -15'd92);
        #4;
        MULT(15'd221, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd126, -15'd19);
        #4;
        MULT(15'd251, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd219, 15'd55);
        #4;
        MULT(15'd77, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd240, 15'd105);
        #4;
        MULT(15'd166, 15'd169);
        #4;
        MULT(15'd35, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd182, -15'd38);
        #4;
        MULT(15'd57, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd17221);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd19, -15'd120);
        #4;
        MULT(15'd203, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd75, -15'd8);
        #4;
        MULT(15'd221, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd115, -15'd36);
        #4;
        MULT(15'd251, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd219, 15'd55);
        #4;
        MULT(15'd77, 15'd55);
        #4;
        MULT(15'd1, 15'd19);
        #4;
        MULT(15'd240, 15'd60);
        #4;
        MULT(15'd166, 15'd105);
        #4;
        MULT(15'd35, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd57, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-76277);
        #4;
        MULT(15'd19, -15'd36);
        #4;
        MULT(15'd203, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd221, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd115, -15'd61);
        #4;
        MULT(15'd52, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd219, 15'd7);
        #4;
        MULT(15'd77, 15'd55);
        #4;
        MULT(15'd1, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd166, 15'd60);
        #4;
        MULT(15'd35, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-134097);
        #4;
        MULT(15'd203, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd115, -15'd100);
        #4;
        MULT(15'd52, -15'd61);
        #4;
        MULT(15'd52, -15'd36);
        #4;
        MULT(15'd219, -15'd19);
        #4;
        MULT(15'd77, 15'd7);
        #4;
        MULT(15'd1, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd35, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-145461);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd219, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd115, -15'd92);
        #4;
        MULT(15'd52, -15'd100);
        #4;
        MULT(15'd52, -15'd61);
        #4;
        MULT(15'd40, -15'd36);
        #4;
        MULT(15'd77, -15'd19);
        #4;
        MULT(15'd1, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-124056);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd219, -15'd3);
        #4;
        MULT(15'd18, -15'd106);
        #4;
        MULT(15'd115, -15'd8);
        #4;
        MULT(15'd52, -15'd92);
        #4;
        MULT(15'd52, -15'd100);
        #4;
        MULT(15'd40, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd1, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-92128);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-4158);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd250, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd229, -15'd82);
        #4;
        CHECK_ACCUM(15'd15186);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd67, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd67, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd250, 15'd197);
        #4;
        MULT(15'd59, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd229, -15'd91);
        #4;
        MULT(15'd21, -15'd82);
        #4;
        CHECK_ACCUM(15'd21276);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd67, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd67, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd250, 15'd169);
        #4;
        MULT(15'd59, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd229, -15'd9);
        #4;
        MULT(15'd21, -15'd91);
        #4;
        MULT(15'd83, -15'd82);
        #4;
        CHECK_ACCUM(15'd-5118);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd67, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd67, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd67, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd250, 15'd105);
        #4;
        MULT(15'd59, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd22, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd229, 15'd102);
        #4;
        MULT(15'd21, -15'd9);
        #4;
        MULT(15'd83, -15'd91);
        #4;
        MULT(15'd233, -15'd82);
        #4;
        CHECK_ACCUM(15'd-36072);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd67, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd67, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd67, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd250, 15'd60);
        #4;
        MULT(15'd59, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd22, 15'd197);
        #4;
        MULT(15'd129, 15'd184);
        #4;
        MULT(15'd229, -15'd38);
        #4;
        MULT(15'd21, 15'd102);
        #4;
        MULT(15'd83, -15'd9);
        #4;
        MULT(15'd233, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd-29810);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd67, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd67, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd59, 15'd19);
        #4;
        MULT(15'd59, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd22, 15'd169);
        #4;
        MULT(15'd129, 15'd197);
        #4;
        MULT(15'd249, 15'd184);
        #4;
        MULT(15'd21, -15'd38);
        #4;
        MULT(15'd83, 15'd102);
        #4;
        MULT(15'd233, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd37016);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd59, 15'd55);
        #4;
        MULT(15'd133, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd22, 15'd105);
        #4;
        MULT(15'd129, 15'd169);
        #4;
        MULT(15'd249, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd83, -15'd38);
        #4;
        MULT(15'd233, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd187, -15'd82);
        #4;
        CHECK_ACCUM(15'd105550);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd9, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd59, 15'd55);
        #4;
        MULT(15'd133, 15'd55);
        #4;
        MULT(15'd205, 15'd19);
        #4;
        MULT(15'd22, 15'd60);
        #4;
        MULT(15'd129, 15'd105);
        #4;
        MULT(15'd249, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd248, 15'd184);
        #4;
        MULT(15'd233, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd187, -15'd91);
        #4;
        MULT(15'd58, -15'd82);
        #4;
        CHECK_ACCUM(15'd159742);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd9, -15'd61);
        #4;
        MULT(15'd126, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd59, 15'd7);
        #4;
        MULT(15'd133, 15'd55);
        #4;
        MULT(15'd205, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd129, 15'd60);
        #4;
        MULT(15'd249, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd248, 15'd197);
        #4;
        MULT(15'd182, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd187, -15'd9);
        #4;
        MULT(15'd58, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd187194);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd75, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd9, -15'd100);
        #4;
        MULT(15'd126, -15'd61);
        #4;
        MULT(15'd251, -15'd36);
        #4;
        MULT(15'd59, -15'd19);
        #4;
        MULT(15'd133, 15'd7);
        #4;
        MULT(15'd205, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd240, 15'd19);
        #4;
        MULT(15'd249, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd248, 15'd169);
        #4;
        MULT(15'd182, 15'd197);
        #4;
        MULT(15'd57, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd187, 15'd102);
        #4;
        MULT(15'd58, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd142807);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd75, -15'd3);
        #4;
        MULT(15'd221, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd9, -15'd92);
        #4;
        MULT(15'd126, -15'd100);
        #4;
        MULT(15'd251, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd133, -15'd19);
        #4;
        MULT(15'd205, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd240, 15'd55);
        #4;
        MULT(15'd166, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd248, 15'd105);
        #4;
        MULT(15'd182, 15'd169);
        #4;
        MULT(15'd57, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd187, -15'd38);
        #4;
        MULT(15'd58, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd49775);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd75, -15'd144);
        #4;
        MULT(15'd221, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd9, -15'd8);
        #4;
        MULT(15'd126, -15'd92);
        #4;
        MULT(15'd251, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd219, -15'd36);
        #4;
        MULT(15'd205, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd240, 15'd55);
        #4;
        MULT(15'd166, 15'd55);
        #4;
        MULT(15'd35, 15'd19);
        #4;
        MULT(15'd248, 15'd60);
        #4;
        MULT(15'd182, 15'd105);
        #4;
        MULT(15'd57, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd58, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-36232);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd75, -15'd120);
        #4;
        MULT(15'd221, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd126, -15'd8);
        #4;
        MULT(15'd251, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd219, -15'd61);
        #4;
        MULT(15'd77, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd240, 15'd7);
        #4;
        MULT(15'd166, 15'd55);
        #4;
        MULT(15'd35, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd182, 15'd60);
        #4;
        MULT(15'd57, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-109327);
        #4;
        MULT(15'd75, -15'd36);
        #4;
        MULT(15'd221, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd115, -15'd106);
        #4;
        MULT(15'd251, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd219, -15'd100);
        #4;
        MULT(15'd77, -15'd61);
        #4;
        MULT(15'd1, -15'd36);
        #4;
        MULT(15'd240, -15'd19);
        #4;
        MULT(15'd166, 15'd7);
        #4;
        MULT(15'd35, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd57, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-128810);
        #4;
        MULT(15'd221, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd115, -15'd3);
        #4;
        MULT(15'd52, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd219, -15'd92);
        #4;
        MULT(15'd77, -15'd100);
        #4;
        MULT(15'd1, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd166, -15'd19);
        #4;
        MULT(15'd35, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-113719);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd115, -15'd144);
        #4;
        MULT(15'd52, -15'd3);
        #4;
        MULT(15'd52, -15'd106);
        #4;
        MULT(15'd219, -15'd8);
        #4;
        MULT(15'd77, -15'd92);
        #4;
        MULT(15'd1, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd35, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-71453);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd115, -15'd120);
        #4;
        MULT(15'd52, -15'd144);
        #4;
        MULT(15'd52, -15'd3);
        #4;
        MULT(15'd40, -15'd106);
        #4;
        MULT(15'd77, -15'd8);
        #4;
        MULT(15'd1, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-35536);
        #4;
        MULT(15'd115, -15'd36);
        #4;
        MULT(15'd52, -15'd120);
        #4;
        MULT(15'd52, -15'd144);
        #4;
        MULT(15'd40, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd1, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-17996);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd198, -15'd82);
        #4;
        CHECK_ACCUM(15'd-4158);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd250, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd229, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd198, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd9196);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd67, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd250, 15'd55);
        #4;
        MULT(15'd59, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd229, 15'd197);
        #4;
        MULT(15'd21, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd198, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd236, -15'd82);
        #4;
        CHECK_ACCUM(15'd-10130);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd67, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd67, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd250, 15'd55);
        #4;
        MULT(15'd59, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd229, 15'd169);
        #4;
        MULT(15'd21, 15'd197);
        #4;
        MULT(15'd83, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd198, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd236, -15'd91);
        #4;
        MULT(15'd253, -15'd82);
        #4;
        CHECK_ACCUM(15'd-35271);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd67, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd67, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd250, 15'd7);
        #4;
        MULT(15'd59, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd22, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd229, 15'd105);
        #4;
        MULT(15'd21, 15'd169);
        #4;
        MULT(15'd83, 15'd197);
        #4;
        MULT(15'd233, 15'd184);
        #4;
        MULT(15'd198, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd236, -15'd9);
        #4;
        MULT(15'd253, -15'd91);
        #4;
        MULT(15'd255, -15'd82);
        #4;
        CHECK_ACCUM(15'd-6233);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd67, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd67, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd250, -15'd19);
        #4;
        MULT(15'd59, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd22, 15'd55);
        #4;
        MULT(15'd129, 15'd19);
        #4;
        MULT(15'd229, 15'd60);
        #4;
        MULT(15'd21, 15'd105);
        #4;
        MULT(15'd83, 15'd169);
        #4;
        MULT(15'd233, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd236, 15'd102);
        #4;
        MULT(15'd253, -15'd9);
        #4;
        MULT(15'd255, -15'd91);
        #4;
        MULT(15'd238, -15'd82);
        #4;
        CHECK_ACCUM(15'd65975);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd67, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd59, -15'd36);
        #4;
        MULT(15'd59, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd22, 15'd55);
        #4;
        MULT(15'd129, 15'd55);
        #4;
        MULT(15'd249, 15'd19);
        #4;
        MULT(15'd21, 15'd60);
        #4;
        MULT(15'd83, 15'd105);
        #4;
        MULT(15'd233, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd236, -15'd38);
        #4;
        MULT(15'd253, 15'd102);
        #4;
        MULT(15'd255, -15'd9);
        #4;
        MULT(15'd238, -15'd91);
        #4;
        MULT(15'd62, -15'd82);
        #4;
        CHECK_ACCUM(15'd140770);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd59, -15'd61);
        #4;
        MULT(15'd133, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd22, 15'd7);
        #4;
        MULT(15'd129, 15'd55);
        #4;
        MULT(15'd249, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd83, 15'd60);
        #4;
        MULT(15'd233, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd187, 15'd184);
        #4;
        MULT(15'd253, -15'd38);
        #4;
        MULT(15'd255, 15'd102);
        #4;
        MULT(15'd238, -15'd9);
        #4;
        MULT(15'd62, -15'd91);
        #4;
        MULT(15'd5, -15'd82);
        #4;
        CHECK_ACCUM(15'd182402);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd9, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd59, -15'd100);
        #4;
        MULT(15'd133, -15'd61);
        #4;
        MULT(15'd205, -15'd36);
        #4;
        MULT(15'd22, -15'd19);
        #4;
        MULT(15'd129, 15'd7);
        #4;
        MULT(15'd249, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd248, 15'd19);
        #4;
        MULT(15'd233, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd187, 15'd197);
        #4;
        MULT(15'd58, 15'd184);
        #4;
        MULT(15'd255, -15'd38);
        #4;
        MULT(15'd238, 15'd102);
        #4;
        MULT(15'd62, -15'd9);
        #4;
        MULT(15'd5, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd155175);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd9, -15'd3);
        #4;
        MULT(15'd126, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd59, -15'd92);
        #4;
        MULT(15'd133, -15'd100);
        #4;
        MULT(15'd205, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd129, -15'd19);
        #4;
        MULT(15'd249, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd248, 15'd55);
        #4;
        MULT(15'd182, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd187, 15'd169);
        #4;
        MULT(15'd58, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd238, -15'd38);
        #4;
        MULT(15'd62, 15'd102);
        #4;
        MULT(15'd5, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd58774);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd9, -15'd144);
        #4;
        MULT(15'd126, -15'd3);
        #4;
        MULT(15'd251, -15'd106);
        #4;
        MULT(15'd59, -15'd8);
        #4;
        MULT(15'd133, -15'd92);
        #4;
        MULT(15'd205, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd240, -15'd36);
        #4;
        MULT(15'd249, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd248, 15'd55);
        #4;
        MULT(15'd182, 15'd55);
        #4;
        MULT(15'd57, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd187, 15'd105);
        #4;
        MULT(15'd58, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd62, -15'd38);
        #4;
        MULT(15'd5, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-21011);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd9, -15'd120);
        #4;
        MULT(15'd126, -15'd144);
        #4;
        MULT(15'd251, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd133, -15'd8);
        #4;
        MULT(15'd205, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd240, -15'd61);
        #4;
        MULT(15'd166, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd248, 15'd7);
        #4;
        MULT(15'd182, 15'd55);
        #4;
        MULT(15'd57, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd187, 15'd60);
        #4;
        MULT(15'd58, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd5, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-85666);
        #4;
        MULT(15'd9, -15'd36);
        #4;
        MULT(15'd126, -15'd120);
        #4;
        MULT(15'd251, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd219, -15'd106);
        #4;
        MULT(15'd205, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd240, -15'd100);
        #4;
        MULT(15'd166, -15'd61);
        #4;
        MULT(15'd35, -15'd36);
        #4;
        MULT(15'd248, -15'd19);
        #4;
        MULT(15'd182, 15'd7);
        #4;
        MULT(15'd57, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd58, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-132781);
        #4;
        MULT(15'd126, -15'd36);
        #4;
        MULT(15'd251, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd219, -15'd3);
        #4;
        MULT(15'd77, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd240, -15'd92);
        #4;
        MULT(15'd166, -15'd100);
        #4;
        MULT(15'd35, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd182, -15'd19);
        #4;
        MULT(15'd57, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-125957);
        #4;
        MULT(15'd251, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd219, -15'd144);
        #4;
        MULT(15'd77, -15'd3);
        #4;
        MULT(15'd1, -15'd106);
        #4;
        MULT(15'd240, -15'd8);
        #4;
        MULT(15'd166, -15'd92);
        #4;
        MULT(15'd35, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd57, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-93164);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd219, -15'd120);
        #4;
        MULT(15'd77, -15'd144);
        #4;
        MULT(15'd1, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd166, -15'd8);
        #4;
        MULT(15'd35, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-51063);
        #4;
        MULT(15'd219, -15'd36);
        #4;
        MULT(15'd77, -15'd120);
        #4;
        MULT(15'd1, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd35, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-17548);
        #4;
        MULT(15'd77, -15'd36);
        #4;
        MULT(15'd1, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2892);
        #4;
        MULT(15'd1, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-36);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd198, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd170, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1862);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd250, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd229, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd198, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd170, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd16089);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd67, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd250, -15'd61);
        #4;
        MULT(15'd59, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd229, 15'd55);
        #4;
        MULT(15'd21, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd198, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd236, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd170, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd254, -15'd82);
        #4;
        CHECK_ACCUM(15'd31786);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd67, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd250, -15'd100);
        #4;
        MULT(15'd59, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd229, 15'd55);
        #4;
        MULT(15'd21, 15'd55);
        #4;
        MULT(15'd83, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd198, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd236, 15'd197);
        #4;
        MULT(15'd253, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd170, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd254, -15'd91);
        #4;
        MULT(15'd209, -15'd82);
        #4;
        CHECK_ACCUM(15'd40923);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd67, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd250, -15'd92);
        #4;
        MULT(15'd59, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd22, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd229, 15'd7);
        #4;
        MULT(15'd21, 15'd55);
        #4;
        MULT(15'd83, 15'd55);
        #4;
        MULT(15'd233, 15'd19);
        #4;
        MULT(15'd198, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd236, 15'd169);
        #4;
        MULT(15'd253, 15'd197);
        #4;
        MULT(15'd255, 15'd184);
        #4;
        MULT(15'd170, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd254, -15'd9);
        #4;
        MULT(15'd209, -15'd91);
        #4;
        MULT(15'd83, -15'd82);
        #4;
        CHECK_ACCUM(15'd95988);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd67, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd250, -15'd8);
        #4;
        MULT(15'd59, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd22, -15'd61);
        #4;
        MULT(15'd129, -15'd36);
        #4;
        MULT(15'd229, -15'd19);
        #4;
        MULT(15'd21, 15'd7);
        #4;
        MULT(15'd83, 15'd55);
        #4;
        MULT(15'd233, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd236, 15'd105);
        #4;
        MULT(15'd253, 15'd169);
        #4;
        MULT(15'd255, 15'd197);
        #4;
        MULT(15'd238, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd254, 15'd102);
        #4;
        MULT(15'd209, -15'd9);
        #4;
        MULT(15'd83, -15'd91);
        #4;
        MULT(15'd44, -15'd82);
        #4;
        CHECK_ACCUM(15'd167422);
        #4;
        MULT(15'd67, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd59, -15'd106);
        #4;
        MULT(15'd59, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd22, -15'd100);
        #4;
        MULT(15'd129, -15'd61);
        #4;
        MULT(15'd249, -15'd36);
        #4;
        MULT(15'd21, -15'd19);
        #4;
        MULT(15'd83, 15'd7);
        #4;
        MULT(15'd233, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd236, 15'd60);
        #4;
        MULT(15'd253, 15'd105);
        #4;
        MULT(15'd255, 15'd169);
        #4;
        MULT(15'd238, 15'd197);
        #4;
        MULT(15'd62, 15'd184);
        #4;
        MULT(15'd254, -15'd38);
        #4;
        MULT(15'd209, 15'd102);
        #4;
        MULT(15'd83, -15'd9);
        #4;
        MULT(15'd44, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd152651);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd59, -15'd3);
        #4;
        MULT(15'd133, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd22, -15'd92);
        #4;
        MULT(15'd129, -15'd100);
        #4;
        MULT(15'd249, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd83, -15'd19);
        #4;
        MULT(15'd233, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd187, 15'd19);
        #4;
        MULT(15'd253, 15'd60);
        #4;
        MULT(15'd255, 15'd105);
        #4;
        MULT(15'd238, 15'd169);
        #4;
        MULT(15'd62, 15'd197);
        #4;
        MULT(15'd5, 15'd184);
        #4;
        MULT(15'd209, -15'd38);
        #4;
        MULT(15'd83, 15'd102);
        #4;
        MULT(15'd44, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd73454);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd59, -15'd144);
        #4;
        MULT(15'd133, -15'd3);
        #4;
        MULT(15'd205, -15'd106);
        #4;
        MULT(15'd22, -15'd8);
        #4;
        MULT(15'd129, -15'd92);
        #4;
        MULT(15'd249, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd248, -15'd36);
        #4;
        MULT(15'd233, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd187, 15'd55);
        #4;
        MULT(15'd58, 15'd19);
        #4;
        MULT(15'd255, 15'd60);
        #4;
        MULT(15'd238, 15'd105);
        #4;
        MULT(15'd62, 15'd169);
        #4;
        MULT(15'd5, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd83, -15'd38);
        #4;
        MULT(15'd44, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-16196);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd59, -15'd120);
        #4;
        MULT(15'd133, -15'd144);
        #4;
        MULT(15'd205, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd129, -15'd8);
        #4;
        MULT(15'd249, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd248, -15'd61);
        #4;
        MULT(15'd182, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd187, 15'd55);
        #4;
        MULT(15'd58, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd238, 15'd60);
        #4;
        MULT(15'd62, 15'd105);
        #4;
        MULT(15'd5, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd44, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-94401);
        #4;
        MULT(15'd59, -15'd36);
        #4;
        MULT(15'd133, -15'd120);
        #4;
        MULT(15'd205, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd240, -15'd106);
        #4;
        MULT(15'd249, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd248, -15'd100);
        #4;
        MULT(15'd182, -15'd61);
        #4;
        MULT(15'd57, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd187, 15'd7);
        #4;
        MULT(15'd58, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd62, 15'd60);
        #4;
        MULT(15'd5, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-133202);
        #4;
        MULT(15'd133, -15'd36);
        #4;
        MULT(15'd205, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd240, -15'd3);
        #4;
        MULT(15'd166, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd248, -15'd92);
        #4;
        MULT(15'd182, -15'd100);
        #4;
        MULT(15'd57, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd187, -15'd19);
        #4;
        MULT(15'd58, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd5, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-133652);
        #4;
        MULT(15'd205, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd240, -15'd144);
        #4;
        MULT(15'd166, -15'd3);
        #4;
        MULT(15'd35, -15'd106);
        #4;
        MULT(15'd248, -15'd8);
        #4;
        MULT(15'd182, -15'd92);
        #4;
        MULT(15'd57, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd58, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-102158);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd240, -15'd120);
        #4;
        MULT(15'd166, -15'd144);
        #4;
        MULT(15'd35, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd182, -15'd8);
        #4;
        MULT(15'd57, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-68653);
        #4;
        MULT(15'd240, -15'd36);
        #4;
        MULT(15'd166, -15'd120);
        #4;
        MULT(15'd35, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd57, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-34056);
        #4;
        MULT(15'd166, -15'd36);
        #4;
        MULT(15'd35, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-10176);
        #4;
        MULT(15'd35, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1260);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd170, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd52, -15'd82);
        #4;
        CHECK_ACCUM(15'd2662);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd250, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd229, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd170, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd52, -15'd91);
        #4;
        MULT(15'd140, -15'd82);
        #4;
        CHECK_ACCUM(15'd32314);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd250, -15'd3);
        #4;
        MULT(15'd59, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd229, -15'd61);
        #4;
        MULT(15'd21, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd198, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd236, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd170, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd254, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd52, -15'd9);
        #4;
        MULT(15'd140, -15'd91);
        #4;
        MULT(15'd106, -15'd82);
        #4;
        CHECK_ACCUM(15'd62907);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd250, -15'd144);
        #4;
        MULT(15'd59, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd229, -15'd100);
        #4;
        MULT(15'd21, -15'd61);
        #4;
        MULT(15'd83, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd198, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd236, 15'd55);
        #4;
        MULT(15'd253, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd170, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd254, 15'd197);
        #4;
        MULT(15'd209, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd52, 15'd102);
        #4;
        MULT(15'd140, -15'd9);
        #4;
        MULT(15'd106, -15'd91);
        #4;
        MULT(15'd18, -15'd82);
        #4;
        CHECK_ACCUM(15'd70013);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd250, -15'd120);
        #4;
        MULT(15'd59, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd22, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd229, -15'd92);
        #4;
        MULT(15'd21, -15'd100);
        #4;
        MULT(15'd83, -15'd61);
        #4;
        MULT(15'd233, -15'd36);
        #4;
        MULT(15'd198, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd236, 15'd55);
        #4;
        MULT(15'd253, 15'd55);
        #4;
        MULT(15'd255, 15'd19);
        #4;
        MULT(15'd170, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd254, 15'd169);
        #4;
        MULT(15'd209, 15'd197);
        #4;
        MULT(15'd83, 15'd184);
        #4;
        MULT(15'd52, -15'd38);
        #4;
        MULT(15'd140, 15'd102);
        #4;
        MULT(15'd106, -15'd9);
        #4;
        MULT(15'd18, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd89550);
        #4;
        MULT(15'd250, -15'd36);
        #4;
        MULT(15'd59, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd22, -15'd3);
        #4;
        MULT(15'd129, -15'd106);
        #4;
        MULT(15'd229, -15'd8);
        #4;
        MULT(15'd21, -15'd92);
        #4;
        MULT(15'd83, -15'd100);
        #4;
        MULT(15'd233, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd236, 15'd7);
        #4;
        MULT(15'd253, 15'd55);
        #4;
        MULT(15'd255, 15'd55);
        #4;
        MULT(15'd238, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd254, 15'd105);
        #4;
        MULT(15'd209, 15'd169);
        #4;
        MULT(15'd83, 15'd197);
        #4;
        MULT(15'd44, 15'd184);
        #4;
        MULT(15'd140, -15'd38);
        #4;
        MULT(15'd106, 15'd102);
        #4;
        MULT(15'd18, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd71055);
        #4;
        MULT(15'd59, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd22, -15'd144);
        #4;
        MULT(15'd129, -15'd3);
        #4;
        MULT(15'd249, -15'd106);
        #4;
        MULT(15'd21, -15'd8);
        #4;
        MULT(15'd83, -15'd92);
        #4;
        MULT(15'd233, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd236, -15'd19);
        #4;
        MULT(15'd253, 15'd7);
        #4;
        MULT(15'd255, 15'd55);
        #4;
        MULT(15'd238, 15'd55);
        #4;
        MULT(15'd62, 15'd19);
        #4;
        MULT(15'd254, 15'd60);
        #4;
        MULT(15'd209, 15'd105);
        #4;
        MULT(15'd83, 15'd169);
        #4;
        MULT(15'd44, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd106, -15'd38);
        #4;
        MULT(15'd18, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-4547);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd22, -15'd120);
        #4;
        MULT(15'd129, -15'd144);
        #4;
        MULT(15'd249, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd83, -15'd8);
        #4;
        MULT(15'd233, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd187, -15'd36);
        #4;
        MULT(15'd253, -15'd19);
        #4;
        MULT(15'd255, 15'd7);
        #4;
        MULT(15'd238, 15'd55);
        #4;
        MULT(15'd62, 15'd55);
        #4;
        MULT(15'd5, 15'd19);
        #4;
        MULT(15'd209, 15'd60);
        #4;
        MULT(15'd83, 15'd105);
        #4;
        MULT(15'd44, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd18, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-77033);
        #4;
        MULT(15'd22, -15'd36);
        #4;
        MULT(15'd129, -15'd120);
        #4;
        MULT(15'd249, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd248, -15'd106);
        #4;
        MULT(15'd233, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd187, -15'd61);
        #4;
        MULT(15'd58, -15'd36);
        #4;
        MULT(15'd255, -15'd19);
        #4;
        MULT(15'd238, 15'd7);
        #4;
        MULT(15'd62, 15'd55);
        #4;
        MULT(15'd5, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd83, 15'd60);
        #4;
        MULT(15'd44, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-133199);
        #4;
        MULT(15'd129, -15'd36);
        #4;
        MULT(15'd249, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd248, -15'd3);
        #4;
        MULT(15'd182, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd187, -15'd100);
        #4;
        MULT(15'd58, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd238, -15'd19);
        #4;
        MULT(15'd62, 15'd7);
        #4;
        MULT(15'd5, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd44, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-139947);
        #4;
        MULT(15'd249, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd248, -15'd144);
        #4;
        MULT(15'd182, -15'd3);
        #4;
        MULT(15'd57, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd187, -15'd92);
        #4;
        MULT(15'd58, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd62, -15'd19);
        #4;
        MULT(15'd5, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-107923);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd248, -15'd120);
        #4;
        MULT(15'd182, -15'd144);
        #4;
        MULT(15'd57, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd187, -15'd8);
        #4;
        MULT(15'd58, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd5, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-72210);
        #4;
        MULT(15'd248, -15'd36);
        #4;
        MULT(15'd182, -15'd120);
        #4;
        MULT(15'd57, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd58, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-39440);
        #4;
        MULT(15'd182, -15'd36);
        #4;
        MULT(15'd57, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-13392);
        #4;
        MULT(15'd57, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2052);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd170, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd52, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-15318);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd229, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd198, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd170, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd52, 15'd197);
        #4;
        MULT(15'd140, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd4090);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd229, -15'd3);
        #4;
        MULT(15'd21, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd198, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd236, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd170, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd52, 15'd169);
        #4;
        MULT(15'd140, 15'd197);
        #4;
        MULT(15'd106, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd8803);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd229, -15'd144);
        #4;
        MULT(15'd21, -15'd3);
        #4;
        MULT(15'd83, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd198, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd236, -15'd61);
        #4;
        MULT(15'd253, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd170, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd209, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd52, 15'd105);
        #4;
        MULT(15'd140, 15'd169);
        #4;
        MULT(15'd106, 15'd197);
        #4;
        MULT(15'd18, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-46302);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd229, -15'd120);
        #4;
        MULT(15'd21, -15'd144);
        #4;
        MULT(15'd83, -15'd3);
        #4;
        MULT(15'd233, -15'd106);
        #4;
        MULT(15'd198, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd236, -15'd100);
        #4;
        MULT(15'd253, -15'd61);
        #4;
        MULT(15'd255, -15'd36);
        #4;
        MULT(15'd170, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd254, 15'd55);
        #4;
        MULT(15'd209, 15'd55);
        #4;
        MULT(15'd83, 15'd19);
        #4;
        MULT(15'd52, 15'd60);
        #4;
        MULT(15'd140, 15'd105);
        #4;
        MULT(15'd106, 15'd169);
        #4;
        MULT(15'd18, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-70874);
        #4;
        MULT(15'd229, -15'd36);
        #4;
        MULT(15'd21, -15'd120);
        #4;
        MULT(15'd83, -15'd144);
        #4;
        MULT(15'd233, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd236, -15'd92);
        #4;
        MULT(15'd253, -15'd100);
        #4;
        MULT(15'd255, -15'd61);
        #4;
        MULT(15'd238, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd254, 15'd7);
        #4;
        MULT(15'd209, 15'd55);
        #4;
        MULT(15'd83, 15'd55);
        #4;
        MULT(15'd44, 15'd19);
        #4;
        MULT(15'd140, 15'd60);
        #4;
        MULT(15'd106, 15'd105);
        #4;
        MULT(15'd18, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-87086);
        #4;
        MULT(15'd21, -15'd36);
        #4;
        MULT(15'd83, -15'd120);
        #4;
        MULT(15'd233, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd236, -15'd8);
        #4;
        MULT(15'd253, -15'd92);
        #4;
        MULT(15'd255, -15'd100);
        #4;
        MULT(15'd238, -15'd61);
        #4;
        MULT(15'd62, -15'd36);
        #4;
        MULT(15'd254, -15'd19);
        #4;
        MULT(15'd209, 15'd7);
        #4;
        MULT(15'd83, 15'd55);
        #4;
        MULT(15'd44, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd106, 15'd60);
        #4;
        MULT(15'd18, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-127496);
        #4;
        MULT(15'd83, -15'd36);
        #4;
        MULT(15'd233, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd187, -15'd106);
        #4;
        MULT(15'd253, -15'd8);
        #4;
        MULT(15'd255, -15'd92);
        #4;
        MULT(15'd238, -15'd100);
        #4;
        MULT(15'd62, -15'd61);
        #4;
        MULT(15'd5, -15'd36);
        #4;
        MULT(15'd209, -15'd19);
        #4;
        MULT(15'd83, 15'd7);
        #4;
        MULT(15'd44, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd18, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-141244);
        #4;
        MULT(15'd233, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd187, -15'd3);
        #4;
        MULT(15'd58, -15'd106);
        #4;
        MULT(15'd255, -15'd8);
        #4;
        MULT(15'd238, -15'd92);
        #4;
        MULT(15'd62, -15'd100);
        #4;
        MULT(15'd5, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd83, -15'd19);
        #4;
        MULT(15'd44, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-113863);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd187, -15'd144);
        #4;
        MULT(15'd58, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd238, -15'd8);
        #4;
        MULT(15'd62, -15'd92);
        #4;
        MULT(15'd5, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd44, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-75670);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd187, -15'd120);
        #4;
        MULT(15'd58, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd62, -15'd8);
        #4;
        MULT(15'd5, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-40892);
        #4;
        MULT(15'd187, -15'd36);
        #4;
        MULT(15'd58, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd5, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-13732);
        #4;
        MULT(15'd58, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2088);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd198, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd170, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd52, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-26120);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd198, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd170, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd52, 15'd55);
        #4;
        MULT(15'd140, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-41512);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd198, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd236, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd170, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd52, 15'd55);
        #4;
        MULT(15'd140, 15'd55);
        #4;
        MULT(15'd106, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-83354);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd198, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd236, -15'd3);
        #4;
        MULT(15'd253, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd170, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd254, -15'd61);
        #4;
        MULT(15'd209, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd52, 15'd7);
        #4;
        MULT(15'd140, 15'd55);
        #4;
        MULT(15'd106, 15'd55);
        #4;
        MULT(15'd18, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-137684);
        #4;
        MULT(15'd198, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd236, -15'd144);
        #4;
        MULT(15'd253, -15'd3);
        #4;
        MULT(15'd255, -15'd106);
        #4;
        MULT(15'd170, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd254, -15'd100);
        #4;
        MULT(15'd209, -15'd61);
        #4;
        MULT(15'd83, -15'd36);
        #4;
        MULT(15'd52, -15'd19);
        #4;
        MULT(15'd140, 15'd7);
        #4;
        MULT(15'd106, 15'd55);
        #4;
        MULT(15'd18, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-158434);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd236, -15'd120);
        #4;
        MULT(15'd253, -15'd144);
        #4;
        MULT(15'd255, -15'd3);
        #4;
        MULT(15'd238, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd254, -15'd92);
        #4;
        MULT(15'd209, -15'd100);
        #4;
        MULT(15'd83, -15'd61);
        #4;
        MULT(15'd44, -15'd36);
        #4;
        MULT(15'd140, -15'd19);
        #4;
        MULT(15'd106, 15'd7);
        #4;
        MULT(15'd18, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-153764);
        #4;
        MULT(15'd236, -15'd36);
        #4;
        MULT(15'd253, -15'd120);
        #4;
        MULT(15'd255, -15'd144);
        #4;
        MULT(15'd238, -15'd3);
        #4;
        MULT(15'd62, -15'd106);
        #4;
        MULT(15'd254, -15'd8);
        #4;
        MULT(15'd209, -15'd92);
        #4;
        MULT(15'd83, -15'd100);
        #4;
        MULT(15'd44, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd106, -15'd19);
        #4;
        MULT(15'd18, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-116994);
        #4;
        MULT(15'd253, -15'd36);
        #4;
        MULT(15'd255, -15'd120);
        #4;
        MULT(15'd238, -15'd144);
        #4;
        MULT(15'd62, -15'd3);
        #4;
        MULT(15'd5, -15'd106);
        #4;
        MULT(15'd209, -15'd8);
        #4;
        MULT(15'd83, -15'd92);
        #4;
        MULT(15'd44, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd18, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-88746);
        #4;
        MULT(15'd255, -15'd36);
        #4;
        MULT(15'd238, -15'd120);
        #4;
        MULT(15'd62, -15'd144);
        #4;
        MULT(15'd5, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd83, -15'd8);
        #4;
        MULT(15'd44, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-51395);
        #4;
        MULT(15'd238, -15'd36);
        #4;
        MULT(15'd62, -15'd120);
        #4;
        MULT(15'd5, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd44, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-17080);
        #4;
        MULT(15'd62, -15'd36);
        #4;
        MULT(15'd5, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-2832);
        #4;
        MULT(15'd5, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-180);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd170, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd52, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-19892);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd170, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd52, -15'd61);
        #4;
        MULT(15'd140, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-35646);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd170, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd254, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd52, -15'd100);
        #4;
        MULT(15'd140, -15'd61);
        #4;
        MULT(15'd106, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-69722);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd170, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd254, -15'd3);
        #4;
        MULT(15'd209, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd52, -15'd92);
        #4;
        MULT(15'd140, -15'd100);
        #4;
        MULT(15'd106, -15'd61);
        #4;
        MULT(15'd18, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-105790);
        #4;
        MULT(15'd170, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd254, -15'd144);
        #4;
        MULT(15'd209, -15'd3);
        #4;
        MULT(15'd83, -15'd106);
        #4;
        MULT(15'd52, -15'd8);
        #4;
        MULT(15'd140, -15'd92);
        #4;
        MULT(15'd106, -15'd100);
        #4;
        MULT(15'd18, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-107595);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd254, -15'd120);
        #4;
        MULT(15'd209, -15'd144);
        #4;
        MULT(15'd83, -15'd3);
        #4;
        MULT(15'd44, -15'd106);
        #4;
        MULT(15'd140, -15'd8);
        #4;
        MULT(15'd106, -15'd92);
        #4;
        MULT(15'd18, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-87305);
        #4;
        MULT(15'd254, -15'd36);
        #4;
        MULT(15'd209, -15'd120);
        #4;
        MULT(15'd83, -15'd144);
        #4;
        MULT(15'd44, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd106, -15'd8);
        #4;
        MULT(15'd18, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-48812);
        #4;
        MULT(15'd209, -15'd36);
        #4;
        MULT(15'd83, -15'd120);
        #4;
        MULT(15'd44, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd18, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-23964);
        #4;
        MULT(15'd83, -15'd36);
        #4;
        MULT(15'd44, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-8268);
        #4;
        MULT(15'd44, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-1584);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd52, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-5512);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd52, -15'd3);
        #4;
        MULT(15'd140, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-14996);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd52, -15'd144);
        #4;
        MULT(15'd140, -15'd3);
        #4;
        MULT(15'd106, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-19144);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd52, -15'd120);
        #4;
        MULT(15'd140, -15'd144);
        #4;
        MULT(15'd106, -15'd3);
        #4;
        MULT(15'd18, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-28626);
        #4;
        MULT(15'd52, -15'd36);
        #4;
        MULT(15'd140, -15'd120);
        #4;
        MULT(15'd106, -15'd144);
        #4;
        MULT(15'd18, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-33990);
        #4;
        MULT(15'd140, -15'd36);
        #4;
        MULT(15'd106, -15'd120);
        #4;
        MULT(15'd18, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-20352);
        #4;
        MULT(15'd106, -15'd36);
        #4;
        MULT(15'd18, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-5976);
        #4;
        MULT(15'd18, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd-648);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd120);
        #4;
        MULT(15'd0, -15'd144);
        #4;
        MULT(15'd0, -15'd3);
        #4;
        MULT(15'd0, -15'd106);
        #4;
        MULT(15'd0, -15'd8);
        #4;
        MULT(15'd0, -15'd92);
        #4;
        MULT(15'd0, -15'd100);
        #4;
        MULT(15'd0, -15'd61);
        #4;
        MULT(15'd0, -15'd36);
        #4;
        MULT(15'd0, -15'd19);
        #4;
        MULT(15'd0, 15'd7);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd55);
        #4;
        MULT(15'd0, 15'd19);
        #4;
        MULT(15'd0, 15'd60);
        #4;
        MULT(15'd0, 15'd105);
        #4;
        MULT(15'd0, 15'd169);
        #4;
        MULT(15'd0, 15'd197);
        #4;
        MULT(15'd0, 15'd184);
        #4;
        MULT(15'd0, -15'd38);
        #4;
        MULT(15'd0, 15'd102);
        #4;
        MULT(15'd0, -15'd9);
        #4;
        MULT(15'd0, -15'd91);
        #4;
        MULT(15'd0, -15'd82);
        #4;
        CHECK_ACCUM(15'd0);

        
        $display("Simulation finished with %d errors", error_count);
				$stop;
        
      end
  
  // Task to simulate key press
  task MULT ( input [15:0] data_fed, input [15:0] weight_fed );
		begin
			data_in = data_fed;
			weight_in = weight_fed;
        	enable = 1'b1;
        	@ (negedge clock) enable = 1'b0;
		end
	endtask
	
			
// Task to check output
  task CHECK_ACCUM ( input [15:0] expResult );
		begin
          
          if (result !== expResult)
				begin
					error_count = error_count + 1;
				end
          reset = 1'b1;
    	@ (negedge clock);
    	@ (negedge clock) reset = 1'b0;
		end
	endtask
	
      
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(2);
  end
endmodule